`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:29:15 10/20/2022 
// Design Name: 
// Module Name:    switchAndLed 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module switchAndLed(switch, led);

	input [7:0] switch;
	output reg [7:0] led;
	
	always@(*)begin
		led = switch;
	end

endmodule
